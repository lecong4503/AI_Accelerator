`timescale 1ns / 1ps

module cnn_kernel